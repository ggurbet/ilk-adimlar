// Gökhan Gurbetoğlu
// GitHub: https://github.com/ggurbet
// Twitter: https://twitter.com/ggurbet
// Programlama Dili: Verilog

module merhaba_dunya ;

initial begin
  $display ("Merhaba Dünya");
  #10  $finish;
end

endmodule
